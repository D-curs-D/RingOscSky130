magic
tech sky130A
timestamp 1637785295
<< locali >>
rect 0 35 27 45
rect 0 15 5 35
rect 22 15 27 35
rect 1155 33 1182 45
rect 1155 25 1160 33
rect 0 0 27 15
rect 1177 25 1182 33
rect 1177 13 1180 25
<< viali >>
rect 5 15 22 35
rect 1160 13 1177 33
<< metal1 >>
rect 0 469 49 735
rect 0 93 49 359
rect 0 35 27 45
rect 0 15 5 35
rect 22 25 27 35
rect 1155 33 1182 45
rect 1155 25 1160 33
rect 22 15 1160 25
rect 0 13 1160 15
rect 1177 13 1182 33
rect 0 0 1182 13
use inv_1  inv_1_2
timestamp 1637503053
transform 1 0 1017 0 1 76
box -229 -76 165 705
use inv_1  inv_1_1
timestamp 1637503053
transform 1 0 623 0 1 76
box -229 -76 165 705
use inv_1  inv_1_0
timestamp 1637503053
transform 1 0 229 0 1 76
box -229 -76 165 705
<< labels >>
rlabel metal1 1177 0 1182 45 3 Y
port 2 e
rlabel space 0 91 49 361 7 VSS
rlabel space 0 466 49 736 7 VDD
rlabel metal1 0 469 49 735 7 VDD
port 1 w
rlabel metal1 0 93 49 359 7 VSS
port 3 w
rlabel space 0 91 49 361 1 remove
<< end >>
